/*
module test (a, b, c);
input signed wire [7:0] a, b;
output signed wire [8:0] c;





endmodule
*/